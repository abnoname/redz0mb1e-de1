------------------------------------------------------------------------------
-- Project    : Red Zombie
------------------------------------------------------------------------------
-- File       :  video_ram_pkg.vhd
-- Author     :  fpgakuechle
-- Company    :  hobbyist
-- Created    :  2012-12
-- Last update: 2013-03-16
-- Licence    : GNU General Public License (http://www.gnu.de/documents/gpl.de.html)
------------------------------------------------------------------------------
-- Description: 
-- used by video_ram.vhd
-- Video memory
-- types and powerUp screen
------------------------------------------------------------------------------
--Last Change: Init Screen with borders, using hexnumbers in index

library ieee;
use ieee.std_logic_1164.all;

package video_ram_pkg is
  SUBTYPE T_VRAM_INDEX IS integer RANGE  0 TO 2**10 - 1;
  SUBTYPE T_WORD       IS integer RANGE 2**8  - 1 DOWNTO 0;
  TYPE    T_VRAM       IS ARRAY (T_VRAM_INDEX'low TO T_VRAM_INDEX'high) OF T_WORD;

--POWERUP screen as initvalues for videoram
  --character tests: letters and digits
  constant C_VRAM_ARRAY_INIT : T_VRAM := (
    --first line
    16#000# => 16#0BC#, 16#001# to 16#01E# => 16#B6#, 16#01F# => 16#BD#,
    --2nd line: col index
    16#020# => 16#B4#,
    16#021# => 16#31#, 16#022# => 16#32#, 16#023# => 16#33#, 16#024# => 16#34#,
    16#025# => 16#35#, 16#026# => 16#36#, 16#027# => 16#37#, 16#028# => 16#38#,
    16#029# => 16#39#, 16#02A# => 16#30#, 16#02B# => 16#31#, 16#02C# => 16#32#,
    16#02D# => 16#33#, 16#02E# => 16#34#, 16#02F# => 16#35#, 

    16#030# => 16#36#,
    16#031# => 16#37#, 16#032# => 16#38#, 16#033# => 16#39#, 16#034# => 16#30#,
    16#035# => 16#31#, 16#036# => 16#32#, 16#037# => 16#33#, 16#038# => 16#34#,
    16#039# => 16#35#, 16#03A# => 16#36#, 16#03B# => 16#37#, 16#03C# => 16#38#,
    16#03D# => 16#39#, 16#03E# => 16#30#,  
    16#03F# => 16#B5#,

    --2nd line: 0x30 - x3F digits and relation
    --0x40- x4F capital letters
--    42 => 16#40#, 43 => 16#41#, 44 => 16#42#, 45 => 16#43#, 46 => 16#44#, 47 => 16#45#, 48 => 16#46#, 49 => 16#47#,
--    52 => 16#48#, 53 => 16#49#, 54 => 16#4A#, 55 => 16#4B#, 56 => 16#4C#, 57 => 16#4D#, 58 => 16#4E#, 59 => 16#4F#,
    --0x50- x5F capital letters
    74 => 16#50#, 75 => 16#51#, 76 => 16#52#, 77 => 16#53#, 78 => 16#54#, 79 => 16#55#, 80 => 16#56#, 81 => 16#57#,
    84 => 16#58#, 85 => 16#59#, 86 => 16#5A#, 87 => 16#5B#, 88 => 16#5C#, 89 => 16#5D#, 90 => 16#5E#, 91 => 16#5F#,
    --0x60- x6F small letter
    106 => 16#60#, 107 => 16#61#, 108 => 16#62#, 109 => 16#63#, 110 => 16#64#, 111 => 16#65#, 112 => 16#66#, 113 => 16#67#,
    116 => 16#68#, 117 => 16#69#, 118 => 16#6A#, 119 => 16#6B#, 120 => 16#6C#, 121 => 16#6D#, 122 => 16#6E#, 123 => 16#6F#,
    --0x70- x7F small letter
    138 => 16#70#, 139 => 16#71#, 140 => 16#72#, 141 => 16#73#, 142 => 16#74#, 143 => 16#75#, 144 => 16#76#, 145 => 16#77#,
    148 => 16#78#, 149 => 16#79#, 150 => 16#7A#, 151 => 16#7B#, 152 => 16#7C#, 153 => 16#7D#, 154 => 16#7E#, 155 => 16#7F#,
    --last line
    16#3E0#  => 16#BB#, 16#3E1# to 16#3FE# => 16#B7#, 16#3FF# => 16#BA#,

    --left border
    16#040# => 16#B4#, 16#041# => 16#32#,
    16#060# => 16#B4#, 16#061# => 16#33#,
    16#080# => 16#B4#, 16#081# => 16#34#,
    16#0A0# => 16#B4#, 16#0A1# => 16#35#,
    16#0C0# => 16#B4#, 16#0C1# => 16#36#,
    16#0E0# => 16#B4#, 16#0E1# => 16#37#,
    16#100# => 16#B4#, 16#101# => 16#38#,
    16#120# => 16#B4#, 16#121# => 16#39#,
    16#140# => 16#B4#, 16#141# => 16#30#,
    16#160# => 16#B4#, 16#161# => 16#31#,
    16#180# => 16#B4#, 16#181# => 16#32#,
    16#1A0# => 16#B4#, 16#1A1# => 16#33#,
    16#1C0# => 16#B4#, 16#1C1# => 16#34#,
    16#1E0# => 16#B4#, 16#1E1# => 16#35#,
    16#200# => 16#B4#, 16#201# => 16#36#,
    16#220# => 16#B4#, 16#221# => 16#37#,
    16#240# => 16#B4#, 16#241# => 16#38#,
    16#260# => 16#B4#, 16#261# => 16#39#,
    16#280# => 16#B4#, 16#281# => 16#30#,
    16#2A0# => 16#B4#, 16#2A1# => 16#31#,
    16#2C0# => 16#B4#, 16#2C1# => 16#32#,
    16#2E0# => 16#B4#, 16#2E1# => 16#33#,
    16#300# => 16#B4#, 16#301# => 16#34#,
    16#320# => 16#B4#, 16#321# => 16#35#,
    16#340# => 16#B4#, 16#341# => 16#36#,
    16#360# => 16#B4#, 16#361# => 16#37#,
    16#380# => 16#B4#, 16#381# => 16#38#,
    16#3A0# => 16#B4#, 16#3A1# => 16#39#,
    16#3C0# => 16#B4#, 16#3C1# => 16#30#,
    -- right border
    16#05F# => 16#B5#, 16#05E# => 16#32#,
    16#07F# => 16#B5#, 16#07E# => 16#33#,
    16#09F# => 16#B5#, 16#09E# => 16#34#,
    16#0BF# => 16#B5#, 16#0BE# => 16#35#,
    16#0DF# => 16#B5#, 16#0DE# => 16#36#,
    16#0FF# => 16#B5#, 16#0FE# => 16#37#,
    16#11F# => 16#B5#, 16#11E# => 16#38#,
    16#13F# => 16#B5#, 16#13E# => 16#39#,
    16#15F# => 16#B5#, 16#15E# => 16#30#,
    16#17F# => 16#B5#, 16#17E# => 16#31#,
    16#19F# => 16#B5#, 16#19E# => 16#32#,
    16#1BF# => 16#B5#, 16#1BE# => 16#33#,
    16#1DF# => 16#B5#, 16#1DE# => 16#34#,
    16#1FF# => 16#B5#, 16#1FE# => 16#35#,
    16#21F# => 16#B5#, 16#21E# => 16#36#,
    16#23F# => 16#B5#, 16#23E# => 16#37#,
    16#25F# => 16#B5#, 16#25E# => 16#38#,
    16#27F# => 16#B5#, 16#27E# => 16#39#,
    16#29F# => 16#B5#, 16#29E# => 16#30#,
    16#2BF# => 16#B5#, 16#2BE# => 16#31#,
    16#2DF# => 16#B5#, 16#2DE# => 16#32#,
    16#2FF# => 16#B5#, 16#2FE# => 16#33#,
    16#31F# => 16#B5#, 16#31E# => 16#34#,
    16#33F# => 16#B5#, 16#33E# => 16#35#,
    16#35F# => 16#B5#, 16#35E# => 16#36#,
    16#37F# => 16#B5#, 16#37E# => 16#37#,
    16#39F# => 16#B5#, 16#39E# => 16#38#,
    16#3BF# => 16#B5#, 16#3BE# => 16#39#,
    16#3DF# => 16#B5#, 16#3DE# => 16#30#,
    others => 16#20#);
  --only spaces -> blank screen
    constant C_VRAM_ARRAY_SPACES_INIT : T_VRAM := (others => 16#20#);
end package video_ram_pkg;

